// System_tb.v

// Generated using ACDS version 13.0sp1 232 at 2025.12.23.15:33:59

`timescale 1 ps / 1 ps
module System_tb (
	);

	wire    system_inst_clk_bfm_clk_clk;          // System_inst_clk_bfm:clk -> [System_inst:clk_clk, System_inst_dma_debug_wm_done_bfm:clk, System_inst_reset_bfm:clk]
	wire    system_inst_reset_bfm_reset_reset;    // System_inst_reset_bfm:reset -> [System_inst:reset_reset_n, System_inst_dma_debug_wm_done_bfm:reset]
	wire    system_inst_dma_debug_wm_done_export; // System_inst:dma_debug_wm_done_export -> System_inst_dma_debug_wm_done_bfm:sig_export

	System system_inst (
		.clk_clk                  (system_inst_clk_bfm_clk_clk),          //               clk.clk
		.reset_reset_n            (system_inst_reset_bfm_reset_reset),    //             reset.reset_n
		.dma_debug_wm_done_export (system_inst_dma_debug_wm_done_export)  // dma_debug_wm_done.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) system_inst_clk_bfm (
		.clk (system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) system_inst_reset_bfm (
		.reset (system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm system_inst_dma_debug_wm_done_bfm (
		.clk        (system_inst_clk_bfm_clk_clk),          //     clk.clk
		.reset      (~system_inst_reset_bfm_reset_reset),   //   reset.reset
		.sig_export (system_inst_dma_debug_wm_done_export)  // conduit.export
	);

endmodule
