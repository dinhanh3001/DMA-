library verilog;
use verilog.vl_types.all;
entity System_tb is
end System_tb;
