module DMAFinal(iClk, iReset_n, iChipselect_n, iRead, iWrite, iAddress, iWritedata, oReaddata, iRM_readdatavalid, iRM_waitrequest, 
iRM_readdata, oRM_read,  oRM_readaddress, iWM_waitrequest, oWM_write, oWM_writeaddress, oWM_writedata, 
   debug_WM_done);
//control slave
input iClk, iReset_n, iChipselect_n, iRead, iWrite;
input [2:0] iAddress;
input [31:0] iWritedata;

output debug_WM_done;   // THEM TIN HIEU DEBUG (SIGNAL TAG) 
output [31:0] oReaddata;
//read master
input iRM_readdatavalid, iRM_waitrequest;
input [31:0] iRM_readdata;

output oRM_read;
output [31:0] oRM_readaddress; 
//write master
input iWM_waitrequest;
output oWM_write;
output [31:0] oWM_writeaddress, oWM_writedata;

wire [31:0] RM_startaddress, length, WM_startaddress, FF_data, FF_q;
wire start, WM_done, FF_almostfull, FF_writerequest, FF_empty, FF_readrequest;

//module control_slave (iClk, iReset_n, iChipselect_n, iWrite, iRead, iMW_done, iAddress, iWritedata,
//						oStart, oReaddata, oRM_startaddress, oWM_startaddress, oLength);
control_slave control(.iClk(iClk), .iReset_n(iReset_n), .iChipselect_n(iChipselect_n), .iWrite(iWrite), .iRead(iRead), 
								.iMW_done(WM_done), .iAddress(iAddress), .iWritedata(iWritedata), .oStart(start), 
								.oReaddata(oReaddata), .oRM_startaddress(RM_startaddress), .oWM_startaddress(WM_startaddress), .oLength(length));

//module write_master ( iClk, iReset_n, iStart, iWM_startaddress, iLength, iWM_waitrequest, iFF_empty, iFF_q, 
//						oFF_readrequest, oWM_done, oWM_write, oWM_writeaddress, oWM_writedata);

write_master wm( .iClk(iClk), .iReset_n(iReset_n), .iStart(start), .iWM_startaddress(WM_startaddress), .iLength(length), .iWM_waitrequest(iWM_waitrequest), .iFF_empty(FF_empty), 
				.iFF_q(FF_q), .oFF_readrequest(FF_readrequest), .oWM_done(WM_done), .oWM_write(oWM_write), .oWM_writeaddress(oWM_writeaddress), .oWM_writedata(oWM_writedata));

					//module read_master(iClk, iReset_n, iStart, iLength, iRM_startaddress, iRM_readdatavalid, iRM_waitrequest
//					oRM_read, oRM_readaddress, iRM_readdata, iFF_almostfull, oFF_writerequest, oFF_data);

read_master rm(.iClk(iClk), .iReset_n(iReset_n), .iStart(start), .iLength(length), .iRM_startaddress(RM_startaddress), .iRM_readdatavalid(iRM_readdatavalid), .iRM_waitrequest(iRM_waitrequest),
					.oRM_read(oRM_read), .oRM_readaddress(oRM_readaddress), .iRM_readdata(iRM_readdata), .iFF_almostfull(FF_almostfull), .oFF_writerequest(FF_writerequest), .oFF_data(FF_data));

//module FIFO(iClk, iReset_n, FF_empty, FF_almostfull, FF_data, FF_q , FF_readrequest, FF_writerequest);

FIFO fi(.iClk(iClk), .iReset_n(iReset_n), .FF_empty(FF_empty), .FF_almostfull(FF_almostfull), .FF_data(FF_data), .FF_q(FF_q) , .FF_readrequest(FF_readrequest), .FF_writerequest(FF_writerequest));
//module fifo (aclr,	clock,data,	rdreq,	wrreq,	almost_full,	empty,	q);
//fifo fi(.aclr(iReset_n),	.clock(iClk), .data(FF_data),	.rdreq(FF_readrequest),	.wrreq(FF_writerequest),	.almost_full(FF_almostfull),	.empty(FF_empty),	.q(FF_q));

assign debug_WM_done = WM_done; 

endmodule 