library verilog;
use verilog.vl_types.all;
entity System_nios2_qsys_0_nios2_performance_monitors is
end System_nios2_qsys_0_nios2_performance_monitors;
